netcdf file\:/D\:/File_2017/T639_Convert/fr/data/201707070852\.NC {
  dimensions:
    x = 104;
    o = 1;
  variables:
    float LON(x);
      LON:long_name = "Flash Longitude";
      LON:standard_name = "Flash Longitude";
      LON:_Unsigned = "FALSE";
      LON:FillValue = 65535.0f;
      LON:valid_range = -180.0f, 180.0f;
      LON:scale_factor = 1.0f;
      LON:add_offset = 0.0f;
      LON:units = "degree";
      LON:resolution = "7800m";
      LON:coordinates = "x";
      LON:ancillary_variables = "DQF";
      LON:_ChunkSizes = 104;

    float LAT(x);
      LAT:long_name = "Flash Latitude";
      LAT:standard_name = "Flash Latitude";
      LAT:_Unsigned = "FALSE";
      LAT:FillValue = 65535.0f;
      LAT:valid_range = -90.0f, 90.0f;
      LAT:scale_factor = 1.0f;
      LAT:add_offset = 0.0f;
      LAT:units = "degree";
      LAT:resolution = "7800m";
      LAT:coordinates = "x";
      LAT:ancillary_variables = "DQF";
      LAT:_ChunkSizes = 104;

    float FTT(x);
      FTT:long_name = "Flash TAI Time";
      FTT:standard_name = "Flash TAI Time";
      FTT:_Unsigned = "FALSE";
      FTT:FillValue = 0.0f;
      FTT:valid_range = 0.0f, 4.0E9f;
      FTT:scale_factor = 1.0f;
      FTT:add_offset = 0.0f;
      FTT:units = "ms";
      FTT:resolution = "7800m";
      FTT:coordinates = "x";
      FTT:ancillary_variables = "DQF";
      FTT:_ChunkSizes = 104;

    float FDT(x);
      FDT:long_name = "Flash Delta Time";
      FDT:standard_name = "Flash Delta Time";
      FDT:_Unsigned = "FALSE";
      FDT:FillValue = 65535.0f;
      FDT:valid_range = 0.0f, 5000.0f;
      FDT:scale_factor = 1.0f;
      FDT:add_offset = 0.0f;
      FDT:units = "ms";
      FDT:resolution = "7800m";
      FDT:coordinates = "x";
      FDT:ancillary_variables = "DQF";
      FDT:_ChunkSizes = 104;

    float FOT(x);
      FOT:long_name = "Flash Observe Time";
      FOT:standard_name = "Flash Observe Time";
      FOT:_Unsigned = "FALSE";
      FOT:FillValue = 0.0f;
      FOT:valid_range = 0.0f, 4.0E9f;
      FOT:scale_factor = 1.0f;
      FOT:add_offset = 0.0f;
      FOT:units = "ms";
      FOT:resolution = "7800m";
      FOT:coordinates = "x";
      FOT:ancillary_variables = "DQF";
      FOT:_ChunkSizes = 104;

    float FR(x);
      FR:long_name = "Flash Radiance";
      FR:standard_name = "Flash Radiance";
      FR:_Unsigned = "FALSE";
      FR:FillValue = 65535.0f;
      FR:valid_range = 0.0f, 10000.0f;
      FR:scale_factor = 1.0f;
      FR:add_offset = 0.0f;
      FR:units = "??J/m*m/ster";
      FR:resolution = "7800m";
      FR:coordinates = "x";
      FR:ancillary_variables = "DQF";
      FR:_ChunkSizes = 104;

    float FF(x);
      FF:long_name = "Flash Footprint";
      FF:standard_name = "Flash Footprint";
      FF:_Unsigned = "FALSE";
      FF:FillValue = 65535.0f;
      FF:valid_range = 0.0f, 10000.0f;
      FF:scale_factor = 1.0f;
      FF:add_offset = 0.0f;
      FF:units = "km2";
      FF:resolution = "7800m";
      FF:coordinates = "x";
      FF:ancillary_variables = "DQF";
      FF:_ChunkSizes = 104;

    float FA(x);
      FA:long_name = "Flash Address";
      FA:standard_name = "Flash Address";
      FA:_Unsigned = "FALSE";
      FA:FillValue = 4.2949673E9f;
      FA:valid_range = 0.0f, 4.0E9f;
      FA:scale_factor = 1.0f;
      FA:add_offset = 0.0f;
      FA:units = "";
      FA:resolution = "7800m";
      FA:coordinates = "x";
      FA:ancillary_variables = "DQF";
      FA:_ChunkSizes = 104;

    float FGA(x);
      FGA:long_name = "Flash Group Address ";
      FGA:standard_name = "Flash Group Address ";
      FGA:_Unsigned = "FALSE";
      FGA:FillValue = 4.2949673E9f;
      FGA:valid_range = 0.0f, 4.0E9f;
      FGA:scale_factor = 1.0f;
      FGA:add_offset = 0.0f;
      FGA:units = "";
      FGA:resolution = "7800m";
      FGA:coordinates = "x";
      FGA:ancillary_variables = "DQF";
      FGA:_ChunkSizes = 104;

    float FGC(x);
      FGC:long_name = "Flash Group Count";
      FGC:standard_name = "Flash  Group Count";
      FGC:_Unsigned = "FALSE";
      FGC:FillValue = 4.2949673E9f;
      FGC:valid_range = 0.0f, 4.0E9f;
      FGC:scale_factor = 1.0f;
      FGC:add_offset = 0.0f;
      FGC:units = "";
      FGC:resolution = "7800m";
      FGC:coordinates = "x";
      FGC:ancillary_variables = "DQF";
      FGC:_ChunkSizes = 104;

    float FEA(x);
      FEA:long_name = "Flash Event Address ";
      FEA:standard_name = "Flash Event Address ";
      FEA:_Unsigned = "FALSE";
      FEA:FillValue = 4.2949673E9f;
      FEA:valid_range = 0.0f, 4.0E9f;
      FEA:scale_factor = 1.0f;
      FEA:add_offset = 0.0f;
      FEA:units = "";
      FEA:resolution = "7800m";
      FEA:coordinates = "x";
      FEA:ancillary_variables = "DQF";
      FEA:_ChunkSizes = 104;

    byte DQF(x);
      DQF:long_name = "Lightening Flash Data Quality Flag";
      DQF:standard_name = "status_flag";
      DQF:_Unsigned = "FALSE";
      DQF:FillValue = 71B;
      DQF:valid_range = 0B, 0B;
      DQF:units = "";
      DQF:coordinates = "x";
      DQF:flag_values = 0B;
      DQF:flag_meanings = "good_pixel conditionally_usable_pixel out_of_range_pixel no_value_pixel";
      DQF:number_of_qf_values = 0B;
      DQF:_ChunkSizes = 104;

    float nominal_satellite_subpoint_lat(o);
      nominal_satellite_subpoint_lat:long_name = "nominal satellite subpoint latitude (platform latitude)";
      nominal_satellite_subpoint_lat:standard_name = "Latitude";
      nominal_satellite_subpoint_lat:units = "degrees_north";
      nominal_satellite_subpoint_lat:_ChunkSizes = 1;

    float nominal_satellite_subpoint_lon(o);
      nominal_satellite_subpoint_lon:units = "degrees_east";
      nominal_satellite_subpoint_lon:long_name = "nominal satellite subpoint longitude (platformlongitude)";
      nominal_satellite_subpoint_lon:standard_name = "Longitude";
      nominal_satellite_subpoint_lon:_ChunkSizes = 1;

    float nominal_satellite_height(o);
      nominal_satellite_height:units = "km";
      nominal_satellite_height:long_name = "nominal satellite height above GRS 80 ellipsoid(platform altitude)";
      nominal_satellite_height:standard_name = "height_above_reference_ellipsoid";
      nominal_satellite_height:_ChunkSizes = 1;

    float geospatial_lat_lon_extent(o);
      geospatial_lat_lon_extent:long_name = "geospatial latitude and longitude references";
      geospatial_lat_lon_extent:begin_line_number = 0US;
      geospatial_lat_lon_extent:end_line_number = 0US;
      geospatial_lat_lon_extent:begin_pixel_number = 0US;
      geospatial_lat_lon_extent:end_pixel_number = 0US;
      geospatial_lat_lon_extent:RegCenterLat = 0.0f;
      geospatial_lat_lon_extent:RegCentralLon = 0.0f;
      geospatial_lat_lon_extent:RegLength = 0.0f;
      geospatial_lat_lon_extent:RegWidth = 0.0f;
      geospatial_lat_lon_extent:geospatial_lat_units = "degrees_north";
      geospatial_lat_lon_extent:geospatial_lon_units = "degrees_east";
      geospatial_lat_lon_extent:_ChunkSizes = 1;

    int OBIType(o);
      OBIType:OBIType_meanings = "NONE";
      OBIType:long_name = "Observing Type";
      OBIType:standard_name = "OBIType";
      OBIType:OBIType_values = 0, 0, -998653952, -697824;
      OBIType:_ChunkSizes = 1;

    int processing_parm_version_container(o);
      processing_parm_version_container:long_name = "NONE";
      processing_parm_version_container:product_version = "NONE";
      processing_parm_version_container:_ChunkSizes = 1;

    int algorithm_product_version_container(o);
      algorithm_product_version_container:long_name = "container for algorithm package filename and productversionchar* sLongName";
      algorithm_product_version_container:product_version = "NONE";
      algorithm_product_version_container:_ChunkSizes = 1;

  // global attributes:
  :dataset_name = "Lightning Imager One Minute";
  :naming_authority = "NSMC CMA";
  :Institution = "NSMC";
  :Project = "GOES";
  :Conventions = "CF-1.7";
  :Metadata_Conv = "Unidata Dataset Discovery v1.0";
  :standard_name_vocabul = "CF Standard Name Table (v25, 05 July 2013)";
  :Title = "Lightning Imager One Minute";
  :Summary = "";
  :platform_ID = "FY-4A";
  :instrument_type = "FengYun-4A Lightning Imager";
  :instrument_ID = "GEOLI";
  :processing_level = "L2";
  :date_created = "2016-02-01T01:15:20.1Z format is YYYY-MM-DD??T??HH:MM:SS.s??Z??.";
  :production_site = "NSMC";
  :production_environment = "";
  :Version_Of_Software = "V1.0";
  :Software_Revision_Date = "YYYY-MM-DD";
  :scene_id = "Region Disk";
  :spatial_resolution = "7800m at nadir";
  :time_coverage_start = "2016-02-01T01:00:00.1Z format is YYYY-MM-DD??T??HH:MM:SS.s??Z??.";
  :time_coverage_end = "2016-02-01T01:13:20.1Z format is YYYY-MM-DD??T??HH:MM:SS.s??Z??.";
  :Data_Quality = "";
  :L0QualityFlag = "";
  :PosQualityFlag = "";
  :CalQualityFlag = "";
  :PosCorFactor1 = "0";
  :PosCorFactor2 = "0";
 data:
LON =
  {83.99979, 113.79933, 121.69921, 110.89938, 114.24317, 114.299324, 104.69947, 113.79933, 121.09921, 94.69962, 113.699326, 119.09926, 110.80154, 121.69921, 110.59938, 113.599335, 121.29922, 104.69947, 108.11262, 122.4992, 117.99927, 120.69922, 121.70194, 83.79979, 111.09937, 104.22524, 119.19925, 125.29916, 82.438194, 117.59927, 119.59924, 116.99928, 120.299225, 120.69922, 107.89942, 118.899254, 118.599266, 120.89923, 116.899284, 121.69921, 123.09919, 116.99928, 79.99985, 94.99962, 119.57291, 109.89939, 111.599365, 121.70891, 121.399216, 111.79936, 100.89953, 114.99931, 119.36699, 119.34982, 122.5992, 110.89937, 114.59931, 111.09937, 110.999374, 86.19975, 116.69929, 104.19948, 121.76464, 124.699165, 116.1879, 120.49923, 121.399216, 104.71288, 117.59927, 121.399216, 121.69921, 120.41408, 118.199265, 121.62451, 122.39919, 121.499214, 110.79938, 83.399796, 115.30374, 92.69966, 116.79929, 125.872185, 122.099205, 115.9993, 93.31948, 108.399414, 124.58325, 113.99933, 117.59928, 122.2992, 122.099205, 122.099205, 96.599594, 121.19922, 112.99935, 115.908005, 119.19926, 83.0998, 121.399185, 120.599236, 105.99945, 86.099754, 112.49936, 121.69921}
LAT =
  {19.065685, 43.80017, 24.900324, 23.326939, 24.900324, 27.700335, 49.500084, 46.000137, 25.000324, 26.800331, 30.000343, 24.123411, 41.40021, 24.742373, 23.90032, 27.500334, 29.20034, 31.000347, 16.100288, 31.100348, 33.500328, 22.70818, 24.976862, 36.200287, 37.100273, 20.30221, 51.00006, 26.100328, 26.420559, 26.50033, 18.4003, 44.60016, 28.000336, 17.600294, 28.100336, 25.200325, 28.70034, 35.700294, 42.0002, 21.700312, 29.600342, 18.200298, 44.100166, 30.400345, 27.382769, 22.200314, 21.300308, 24.89975, 25.000324, 24.400322, 33.700325, 17.600296, 26.991142, 27.000332, 31.100348, 23.300318, 45.971813, 16.600292, 27.900335, 16.800293, 26.60033, 37.500267, 24.900324, 29.30034, 28.680004, 17.000294, 53.70002, 49.400085, 26.50033, 25.000324, 24.900324, 24.338654, 20.300306, 25.100323, 53.900017, 17.700296, 41.400208, 20.800308, 18.952341, 22.200314, 23.70032, 38.32853, 25.800327, 18.4003, 23.638914, 23.40032, 28.684418, 46.200134, 26.55461, 51.00006, 51.00006, 50.800064, 17.900297, 29.30034, 18.900303, 25.594654, 51.00006, 35.500298, 24.876377, 18.300299, 27.200333, 23.200317, 18.8003, 24.800323}
FTT =
  {240.0, 1500.0, 2600.0, 2978.0, 3782.0, 3920.0, 4072.0, 4392.0, 5010.0, 5932.0, 6324.0, 6840.0, 8230.0, 8238.0, 8298.0, 9682.0, 10096.0, 10856.0, 11764.0, 13224.0, 13722.0, 14784.0, 16346.0, 16460.0, 17094.0, 17614.0, 18240.0, 18364.0, 18534.0, 18936.0, 19446.0, 19466.0, 19584.0, 19974.0, 20204.0, 20534.0, 21686.0, 21768.0, 21972.0, 22244.0, 22964.0, 23014.0, 24020.0, 24208.0, 25374.0, 26564.0, 27268.0, 27394.0, 27432.0, 28656.0, 29092.0, 29758.0, 29866.0, 30314.0, 30706.0, 30736.0, 31388.0, 31544.0, 31748.0, 31872.0, 32308.0, 32364.0, 33258.0, 34170.0, 34210.0, 34486.0, 37502.0, 37864.0, 38202.0, 38302.0, 38404.0, 38418.0, 38824.0, 39602.0, 39748.0, 42994.0, 43332.0, 43692.0, 43878.0, 44016.0, 44082.0, 45288.0, 46236.0, 46502.0, 47328.0, 47352.0, 48532.0, 48592.0, 48636.0, 48864.0, 48864.0, 48864.0, 49562.0, 49676.0, 49820.0, 50246.0, 50500.0, 51218.0, 53010.0, 53458.0, 54592.0, 55512.0, 55690.0, 55796.0}
FDT =
  {2.0, 0.0, 0.0, 0.0, 20.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 90.0, 0.0, 0.0, 0.0, 0.0, 14.0, 0.0, 0.0, 0.0, 222.0, 0.0, 0.0, 18.0, 0.0, 0.0, 2.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 82.0, 30.0, 0.0, 324.0, 0.0, 0.0, 0.0, 0.0, 74.0, 0.0, 0.0, 100.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 72.0, 0.0, 0.0, 0.0, 116.0, 0.0, 0.0, 0.0, 92.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 120.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 218.0, 292.0, 152.0, 0.0, 402.0, 0.0, 0.0, 4.0, 88.0, 0.0}
FOT =
  {100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0}
FR =
  {3.5350397, 3.1816068, 0.7461536, 16.985928, 50.651794, 1.0793892, 2.003521, 4.62065, 2.930124, 1.5981306, 2.8091605, 10.454092, 3.4084928, 12.680096, 3.3471582, 2.6875956, 1.9384613, 0.07283756, 3.345578, 0.40435436, 1.5405406, 6.045507, 13.603853, 2.6119757, 2.1678405, 289.45557, 0.95949084, 0.4901365, 175.83437, 1.1790123, 0.36656433, 4.2587414, 0.38724756, 1.3877778, 1.0531915, 5.265023, 1.4219476, 1.6600466, 2.3528724, 0.44822282, 0.17465241, 4.398723, 20.028402, 4.0833335, 48.34541, 6.6273293, 6.7950306, 45.843502, 2.095827, 0.27469116, 2.73753, 4.426563, 22.095451, 11.649612, 1.306028, 17.121933, 13.039677, 1.5378549, 3.706538, 15.6992, 3.9349468, 3.5475912, 6.608602, 8.365443, 4.84229, 5.611801, 0.09699771, 17.185108, 1.7962962, 0.14660506, 26.247414, 15.259823, 0.24116738, 1.7260484, 3.1020641, 1.848297, 0.056206036, 1.7563692, 43.769234, 124.52602, 3.043546, 52.95334, 0.11230762, 1.6094943, 160.07585, 12.469136, 5.0861516, 4.342625, 13.042278, 159.37798, 139.21844, 3.2760668, 0.6987382, 3.052795, 20.010529, 35.437035, 3.5393517, 2.2422059, 30.031895, 2.9290123, 7.413476, 2.4444435, 6.626521, 1.1843317}
FF =
  {400.0, 100.0, 100.0, 400.0, 700.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 300.0, 200.0, 400.0, 100.0, 100.0, 100.0, 100.0, 300.0, 100.0, 100.0, 200.0, 400.0, 100.0, 100.0, 1800.0, 100.0, 100.0, 1400.0, 100.0, 100.0, 100.0, 100.0, 200.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 200.0, 100.0, 100.0, 900.0, 200.0, 100.0, 700.0, 100.0, 100.0, 100.0, 100.0, 800.0, 200.0, 100.0, 500.0, 200.0, 100.0, 200.0, 100.0, 100.0, 100.0, 200.0, 100.0, 300.0, 100.0, 100.0, 300.0, 100.0, 100.0, 200.0, 700.0, 100.0, 200.0, 100.0, 200.0, 100.0, 100.0, 700.0, 200.0, 100.0, 700.0, 100.0, 100.0, 1000.0, 100.0, 200.0, 100.0, 200.0, 100.0, 100.0, 100.0, 100.0, 100.0, 600.0, 600.0, 200.0, 100.0, 1000.0, 100.0, 100.0, 200.0, 300.0, 100.0}
FA =
  {1.0, 2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0, 46.0, 47.0, 48.0, 49.0, 50.0, 51.0, 52.0, 53.0, 54.0, 55.0, 56.0, 57.0, 58.0, 59.0, 60.0, 61.0, 62.0, 63.0, 64.0, 65.0, 66.0, 67.0, 68.0, 69.0, 70.0, 71.0, 72.0, 73.0, 74.0, 75.0, 76.0, 77.0, 78.0, 79.0, 80.0, 81.0, 82.0, 83.0, 84.0, 85.0, 86.0, 87.0, 88.0, 89.0, 90.0, 91.0, 92.0, 93.0, 94.0, 95.0, 96.0, 97.0, 98.0, 99.0, 100.0, 101.0, 102.0, 103.0, 104.0}
FGA =
  {0.0, 2.0, 3.0, 4.0, 5.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 18.0, 19.0, 20.0, 21.0, 22.0, 24.0, 25.0, 26.0, 27.0, 29.0, 30.0, 31.0, 34.0, 35.0, 36.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0, 46.0, 47.0, 48.0, 49.0, 50.0, 51.0, 52.0, 53.0, 55.0, 57.0, 58.0, 62.0, 63.0, 64.0, 65.0, 66.0, 70.0, 71.0, 72.0, 75.0, 76.0, 77.0, 78.0, 79.0, 80.0, 81.0, 82.0, 83.0, 84.0, 85.0, 86.0, 88.0, 89.0, 90.0, 91.0, 95.0, 96.0, 97.0, 98.0, 100.0, 101.0, 102.0, 103.0, 104.0, 105.0, 106.0, 107.0, 108.0, 111.0, 112.0, 113.0, 114.0, 115.0, 116.0, 117.0, 118.0, 119.0, 120.0, 123.0, 125.0, 127.0, 128.0, 136.0, 137.0, 138.0, 140.0, 142.0}
FGC =
  {2.0, 1.0, 1.0, 1.0, 2.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 3.0, 1.0, 1.0, 1.0, 1.0, 2.0, 1.0, 1.0, 1.0, 2.0, 1.0, 1.0, 3.0, 1.0, 1.0, 2.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 2.0, 2.0, 1.0, 4.0, 1.0, 1.0, 1.0, 1.0, 4.0, 1.0, 1.0, 3.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 2.0, 1.0, 1.0, 1.0, 4.0, 1.0, 1.0, 1.0, 2.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 3.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 3.0, 2.0, 2.0, 1.0, 8.0, 1.0, 1.0, 2.0, 2.0, 1.0}
FEA =
  {4.0, 1.0, 1.0, 4.0, 7.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 3.0, 2.0, 4.0, 1.0, 1.0, 1.0, 1.0, 3.0, 1.0, 1.0, 2.0, 4.0, 1.0, 1.0, 18.0, 1.0, 1.0, 14.0, 1.0, 1.0, 1.0, 1.0, 2.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 2.0, 1.0, 1.0, 9.0, 2.0, 1.0, 7.0, 1.0, 1.0, 1.0, 1.0, 8.0, 2.0, 1.0, 5.0, 2.0, 1.0, 2.0, 1.0, 1.0, 1.0, 2.0, 1.0, 3.0, 1.0, 1.0, 3.0, 1.0, 1.0, 2.0, 7.0, 1.0, 2.0, 1.0, 2.0, 1.0, 1.0, 7.0, 2.0, 1.0, 7.0, 1.0, 1.0, 10.0, 1.0, 2.0, 1.0, 2.0, 1.0, 1.0, 1.0, 1.0, 1.0, 6.0, 6.0, 2.0, 1.0, 10.0, 1.0, 1.0, 2.0, 3.0, 1.0}
DQF =
  {0, 1, 1, 1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 0, 1, 1, 1, 1, 0, 1, 1, 1, 0, 1, 1, 0, 1, 1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 1, 0, 1, 1, 1, 1, 0, 1, 1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 1, 1, 1, 0, 1, 1, 1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 1, 0, 1, 1, 0, 0, 1}
nominal_satellite_subpoint_lat =
  {0.0}
nominal_satellite_subpoint_lon =
  {0.0}
nominal_satellite_height =
  {0.0}
geospatial_lat_lon_extent =
  {0.0}
OBIType =
  {0}
processing_parm_version_container =
  {0}
algorithm_product_version_container =
  {0}
}
