netcdf file\:/D\:/File_2017/T639_Convert/fr/data/201707070851\.NC {
  dimensions:
    x = 109;
    o = 1;
  variables:
    float LON(x);
      LON:long_name = "Flash Longitude";
      LON:standard_name = "Flash Longitude";
      LON:_Unsigned = "FALSE";
      LON:FillValue = 65535.0f;
      LON:valid_range = -180.0f, 180.0f;
      LON:scale_factor = 1.0f;
      LON:add_offset = 0.0f;
      LON:units = "degree";
      LON:resolution = "7800m";
      LON:coordinates = "x";
      LON:ancillary_variables = "DQF";
      LON:_ChunkSizes = 109;

    float LAT(x);
      LAT:long_name = "Flash Latitude";
      LAT:standard_name = "Flash Latitude";
      LAT:_Unsigned = "FALSE";
      LAT:FillValue = 65535.0f;
      LAT:valid_range = -90.0f, 90.0f;
      LAT:scale_factor = 1.0f;
      LAT:add_offset = 0.0f;
      LAT:units = "degree";
      LAT:resolution = "7800m";
      LAT:coordinates = "x";
      LAT:ancillary_variables = "DQF";
      LAT:_ChunkSizes = 109;

    float FTT(x);
      FTT:long_name = "Flash TAI Time";
      FTT:standard_name = "Flash TAI Time";
      FTT:_Unsigned = "FALSE";
      FTT:FillValue = 0.0f;
      FTT:valid_range = 0.0f, 4.0E9f;
      FTT:scale_factor = 1.0f;
      FTT:add_offset = 0.0f;
      FTT:units = "ms";
      FTT:resolution = "7800m";
      FTT:coordinates = "x";
      FTT:ancillary_variables = "DQF";
      FTT:_ChunkSizes = 109;

    float FDT(x);
      FDT:long_name = "Flash Delta Time";
      FDT:standard_name = "Flash Delta Time";
      FDT:_Unsigned = "FALSE";
      FDT:FillValue = 65535.0f;
      FDT:valid_range = 0.0f, 5000.0f;
      FDT:scale_factor = 1.0f;
      FDT:add_offset = 0.0f;
      FDT:units = "ms";
      FDT:resolution = "7800m";
      FDT:coordinates = "x";
      FDT:ancillary_variables = "DQF";
      FDT:_ChunkSizes = 109;

    float FOT(x);
      FOT:long_name = "Flash Observe Time";
      FOT:standard_name = "Flash Observe Time";
      FOT:_Unsigned = "FALSE";
      FOT:FillValue = 0.0f;
      FOT:valid_range = 0.0f, 4.0E9f;
      FOT:scale_factor = 1.0f;
      FOT:add_offset = 0.0f;
      FOT:units = "ms";
      FOT:resolution = "7800m";
      FOT:coordinates = "x";
      FOT:ancillary_variables = "DQF";
      FOT:_ChunkSizes = 109;

    float FR(x);
      FR:long_name = "Flash Radiance";
      FR:standard_name = "Flash Radiance";
      FR:_Unsigned = "FALSE";
      FR:FillValue = 65535.0f;
      FR:valid_range = 0.0f, 10000.0f;
      FR:scale_factor = 1.0f;
      FR:add_offset = 0.0f;
      FR:units = "??J/m*m/ster";
      FR:resolution = "7800m";
      FR:coordinates = "x";
      FR:ancillary_variables = "DQF";
      FR:_ChunkSizes = 109;

    float FF(x);
      FF:long_name = "Flash Footprint";
      FF:standard_name = "Flash Footprint";
      FF:_Unsigned = "FALSE";
      FF:FillValue = 65535.0f;
      FF:valid_range = 0.0f, 10000.0f;
      FF:scale_factor = 1.0f;
      FF:add_offset = 0.0f;
      FF:units = "km2";
      FF:resolution = "7800m";
      FF:coordinates = "x";
      FF:ancillary_variables = "DQF";
      FF:_ChunkSizes = 109;

    float FA(x);
      FA:long_name = "Flash Address";
      FA:standard_name = "Flash Address";
      FA:_Unsigned = "FALSE";
      FA:FillValue = 4.2949673E9f;
      FA:valid_range = 0.0f, 4.0E9f;
      FA:scale_factor = 1.0f;
      FA:add_offset = 0.0f;
      FA:units = "";
      FA:resolution = "7800m";
      FA:coordinates = "x";
      FA:ancillary_variables = "DQF";
      FA:_ChunkSizes = 109;

    float FGA(x);
      FGA:long_name = "Flash Group Address ";
      FGA:standard_name = "Flash Group Address ";
      FGA:_Unsigned = "FALSE";
      FGA:FillValue = 4.2949673E9f;
      FGA:valid_range = 0.0f, 4.0E9f;
      FGA:scale_factor = 1.0f;
      FGA:add_offset = 0.0f;
      FGA:units = "";
      FGA:resolution = "7800m";
      FGA:coordinates = "x";
      FGA:ancillary_variables = "DQF";
      FGA:_ChunkSizes = 109;

    float FGC(x);
      FGC:long_name = "Flash Group Count";
      FGC:standard_name = "Flash  Group Count";
      FGC:_Unsigned = "FALSE";
      FGC:FillValue = 4.2949673E9f;
      FGC:valid_range = 0.0f, 4.0E9f;
      FGC:scale_factor = 1.0f;
      FGC:add_offset = 0.0f;
      FGC:units = "";
      FGC:resolution = "7800m";
      FGC:coordinates = "x";
      FGC:ancillary_variables = "DQF";
      FGC:_ChunkSizes = 109;

    float FEA(x);
      FEA:long_name = "Flash Event Address ";
      FEA:standard_name = "Flash Event Address ";
      FEA:_Unsigned = "FALSE";
      FEA:FillValue = 4.2949673E9f;
      FEA:valid_range = 0.0f, 4.0E9f;
      FEA:scale_factor = 1.0f;
      FEA:add_offset = 0.0f;
      FEA:units = "";
      FEA:resolution = "7800m";
      FEA:coordinates = "x";
      FEA:ancillary_variables = "DQF";
      FEA:_ChunkSizes = 109;

    byte DQF(x);
      DQF:long_name = "Lightening Flash Data Quality Flag";
      DQF:standard_name = "status_flag";
      DQF:_Unsigned = "FALSE";
      DQF:FillValue = 71B;
      DQF:valid_range = 0B, 0B;
      DQF:units = "";
      DQF:coordinates = "x";
      DQF:flag_values = 0B;
      DQF:flag_meanings = "good_pixel conditionally_usable_pixel out_of_range_pixel no_value_pixel";
      DQF:number_of_qf_values = 0B;
      DQF:_ChunkSizes = 109;

    float nominal_satellite_subpoint_lat(o);
      nominal_satellite_subpoint_lat:long_name = "nominal satellite subpoint latitude (platform latitude)";
      nominal_satellite_subpoint_lat:standard_name = "Latitude";
      nominal_satellite_subpoint_lat:units = "degrees_north";
      nominal_satellite_subpoint_lat:_ChunkSizes = 1;

    float nominal_satellite_subpoint_lon(o);
      nominal_satellite_subpoint_lon:units = "degrees_east";
      nominal_satellite_subpoint_lon:long_name = "nominal satellite subpoint longitude (platformlongitude)";
      nominal_satellite_subpoint_lon:standard_name = "Longitude";
      nominal_satellite_subpoint_lon:_ChunkSizes = 1;

    float nominal_satellite_height(o);
      nominal_satellite_height:units = "km";
      nominal_satellite_height:long_name = "nominal satellite height above GRS 80 ellipsoid(platform altitude)";
      nominal_satellite_height:standard_name = "height_above_reference_ellipsoid";
      nominal_satellite_height:_ChunkSizes = 1;

    float geospatial_lat_lon_extent(o);
      geospatial_lat_lon_extent:long_name = "geospatial latitude and longitude references";
      geospatial_lat_lon_extent:begin_line_number = 0US;
      geospatial_lat_lon_extent:end_line_number = 0US;
      geospatial_lat_lon_extent:begin_pixel_number = 0US;
      geospatial_lat_lon_extent:end_pixel_number = 0US;
      geospatial_lat_lon_extent:RegCenterLat = 0.0f;
      geospatial_lat_lon_extent:RegCentralLon = 0.0f;
      geospatial_lat_lon_extent:RegLength = 0.0f;
      geospatial_lat_lon_extent:RegWidth = 0.0f;
      geospatial_lat_lon_extent:geospatial_lat_units = "degrees_north";
      geospatial_lat_lon_extent:geospatial_lon_units = "degrees_east";
      geospatial_lat_lon_extent:_ChunkSizes = 1;

    int OBIType(o);
      OBIType:OBIType_meanings = "NONE";
      OBIType:long_name = "Observing Type";
      OBIType:standard_name = "OBIType";
      OBIType:OBIType_values = 0, 0, -998653952, -697856;
      OBIType:_ChunkSizes = 1;

    int processing_parm_version_container(o);
      processing_parm_version_container:long_name = "NONE";
      processing_parm_version_container:product_version = "NONE";
      processing_parm_version_container:_ChunkSizes = 1;

    int algorithm_product_version_container(o);
      algorithm_product_version_container:long_name = "container for algorithm package filename and productversionchar* sLongName";
      algorithm_product_version_container:product_version = "NONE";
      algorithm_product_version_container:_ChunkSizes = 1;

  // global attributes:
  :dataset_name = "Lightning Imager One Minute";
  :naming_authority = "NSMC CMA";
  :Institution = "NSMC";
  :Project = "GOES";
  :Conventions = "CF-1.7";
  :Metadata_Conv = "Unidata Dataset Discovery v1.0";
  :standard_name_vocabul = "CF Standard Name Table (v25, 05 July 2013)";
  :Title = "Lightning Imager One Minute";
  :Summary = "";
  :platform_ID = "FY-4A";
  :instrument_type = "FengYun-4A Lightning Imager";
  :instrument_ID = "GEOLI";
  :processing_level = "L2";
  :date_created = "2016-02-01T01:15:20.1Z format is YYYY-MM-DD??T??HH:MM:SS.s??Z??.";
  :production_site = "NSMC";
  :production_environment = "";
  :Version_Of_Software = "V1.0";
  :Software_Revision_Date = "YYYY-MM-DD";
  :scene_id = "Region Disk";
  :spatial_resolution = "7800m at nadir";
  :time_coverage_start = "2016-02-01T01:00:00.1Z format is YYYY-MM-DD??T??HH:MM:SS.s??Z??.";
  :time_coverage_end = "2016-02-01T01:13:20.1Z format is YYYY-MM-DD??T??HH:MM:SS.s??Z??.";
  :Data_Quality = "";
  :L0QualityFlag = "";
  :PosQualityFlag = "";
  :CalQualityFlag = "";
  :PosCorFactor1 = "0";
  :PosCorFactor2 = "0";
 data:
LON =
  {111.49936, 119.49925, 113.89933, 113.88713, 106.09945, 108.399414, 94.79962, 109.3994, 120.49014, 84.99977, 115.33795, 123.69917, 108.399414, 105.89945, 114.199326, 133.99948, 133.79947, 116.29929, 117.89927, 119.29925, 105.099464, 87.49973, 99.69955, 117.56987, 98.39957, 121.499214, 98.99956, 113.55146, 121.19922, 116.1993, 128.17007, 121.39535, 120.59923, 115.92309, 92.89965, 113.599335, 113.69933, 121.737854, 114.79932, 114.09933, 125.79915, 108.813644, 114.092606, 96.2996, 83.0998, 110.89938, 119.3777, 92.39966, 102.09951, 109.0994, 116.59929, 92.49966, 127.69913, 123.79918, 112.799355, 104.89947, 101.99951, 121.69921, 104.28926, 118.399254, 108.29941, 110.152695, 115.57709, 111.09937, 119.19925, 106.79944, 125.399155, 118.69926, 86.16541, 105.099464, 125.518654, 119.543976, 123.39919, 121.6992, 125.59915, 117.158844, 117.19928, 111.722115, 84.26067, 119.39925, 97.799576, 118.699265, 88.09293, 118.69926, 108.21702, 114.199326, 87.09974, 117.39928, 87.01848, 86.99974, 121.39922, 107.79942, 113.89436, 110.89168, 110.89938, 114.62584, 112.99935, 98.64438, 121.36043, 121.29922, 115.9758, 108.89941, 120.44115, 120.55104, 111.15932, 119.19925, 118.49926, 123.399185, 94.09963}
LAT =
  {22.689997, 26.900333, 46.100136, 20.35185, 19.400303, 32.200348, 39.700233, 41.600204, 16.918459, 35.90029, 18.95899, 29.957651, 41.700203, 48.600098, 26.800331, 44.800156, 44.800156, 23.700321, 26.70033, 27.000332, 21.20031, 23.300318, 16.900291, 26.518856, 21.800314, 17.800297, 41.700203, 43.652298, 29.30034, 24.10032, 26.300331, 24.999496, 24.432058, 25.584356, 22.600315, 50.800064, 51.00006, 24.897085, 46.000137, 24.900324, 54.600006, 28.700338, 24.900324, 16.900293, 35.500298, 23.30032, 26.931873, 33.600327, 18.300299, 36.800278, 26.30033, 17.200294, 29.800343, 45.10015, 39.700233, 48.5001, 45.30015, 25.000324, 20.290688, 27.396486, 40.800217, 23.01421, 25.571909, 28.000336, 51.00006, 31.300348, 32.10035, 26.60033, 23.164455, 21.20031, 16.500292, 26.800331, 19.600304, 25.100325, 44.100166, 51.995476, 52.200043, 23.904573, 22.155478, 27.000332, 26.100327, 27.00033, 23.269886, 27.000332, 22.90351, 30.600346, 51.80005, 26.500332, 28.681602, 29.10034, 29.400341, 29.800343, 20.276003, 23.402098, 23.30032, 46.000137, 18.900301, 40.41407, 24.946978, 24.743078, 25.582458, 28.700338, 16.858366, 16.943275, 27.897333, 51.00006, 23.80032, 35.100304, 31.70035}
FTT =
  {92.0, 672.0, 1550.0, 2794.0, 4686.0, 5044.0, 5054.0, 5476.0, 6376.0, 6966.0, 7092.0, 7538.0, 7712.0, 7874.0, 8330.0, 8470.0, 8470.0, 8738.0, 8916.0, 8998.0, 9904.0, 10328.0, 10374.0, 10460.0, 11042.0, 11448.0, 11864.0, 12528.0, 13522.0, 13772.0, 13828.0, 16368.0, 16422.0, 16426.0, 16722.0, 17314.0, 17314.0, 17196.0, 17674.0, 17824.0, 18120.0, 18426.0, 18312.0, 19018.0, 19630.0, 20060.0, 21476.0, 21526.0, 21848.0, 22224.0, 25794.0, 26468.0, 26774.0, 26974.0, 27188.0, 27362.0, 27676.0, 28468.0, 28454.0, 28872.0, 31228.0, 31414.0, 32004.0, 32050.0, 32376.0, 32680.0, 33186.0, 33366.0, 33398.0, 33540.0, 33892.0, 35574.0, 35598.0, 35744.0, 36414.0, 38594.0, 38594.0, 39794.0, 39872.0, 40216.0, 40972.0, 40998.0, 41148.0, 41442.0, 41712.0, 43008.0, 43356.0, 44266.0, 44804.0, 44804.0, 44842.0, 45624.0, 45548.0, 45608.0, 47896.0, 48438.0, 49414.0, 49428.0, 49390.0, 50150.0, 50448.0, 50490.0, 51414.0, 51768.0, 52328.0, 52932.0, 53060.0, 53548.0, 53930.0}
FDT =
  {62.0, 100.0, 0.0, 50.0, 0.0, 0.0, 0.0, 0.0, 170.0, 2.0, 64.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 284.0, 0.0, 0.0, 0.0, 6.0, 2.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 334.0, 0.0, 0.0, 0.0, 0.0, 0.0, 326.0, 0.0, 0.0, 0.0, 4.0, 444.0, 0.0, 0.0, 208.0, 280.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 98.0, 0.0, 0.0, 492.0, 36.0, 0.0, 0.0, 0.0, 0.0, 0.0, 78.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 0.0, 126.0, 160.0, 28.0, 0.0, 80.0, 0.0, 0.0, 406.0, 0.0, 2.0, 0.0, 0.0, 0.0, 0.0, 0.0, 440.0, 516.0, 0.0, 2.0, 0.0, 0.0, 820.0, 48.0, 240.0, 0.0, 24.0, 80.0, 252.0, 12.0, 0.0, 0.0, 0.0}
FOT =
  {100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0}
FR =
  {10.620317, 0.75465846, 0.11475404, 199.92697, 3.545171, 0.47938922, 2.254459, 0.13395998, 133.21654, 25.12067, 141.77132, 48.63463, 4.0861864, 3.9834516, 0.25762174, 57.033096, 0.565574, 1.4429222, 14.94847, 0.84378356, 2.3479624, 0.07679993, 5.1943126, 4.634285, 1.6745285, 2.52093, 10.99881, 5.0483427, 1.189441, 2.9737253, 7.7770987, 43.92226, 6.006462, 35.00317, 0.9795278, 20.799072, 0.1104652, 240.60454, 0.89120376, 3.0668695, 1.1785296, 31.746094, 36.11614, 6.4213834, 7.7577934, 36.104336, 69.4368, 0.5597637, 0.9936104, 2.2681499, 1.0627804, 1.5113639, 3.0430768, 0.16273554, 19.184364, 2.6588511, 0.09735548, 1.6609373, 331.11923, 80.95522, 19.010574, 1289.3401, 15.091152, 0.99231935, 0.2650464, 0.97247714, 1.8052148, 10.193846, 1049.772, 2.3479624, 13.50605, 3.7730613, 1.2083334, 0.28081113, 8.082944, 50.767273, 2.3213036, 14.712872, 249.56561, 3.7209303, 19.997663, 2.9306622, 255.4501, 0.4637902, 281.07544, 0.24542692, 8.012152, 1.2703533, 117.44759, 1.0218071, 4.373272, 6.8088684, 417.5583, 764.8305, 2.7833166, 17.061062, 4.3804574, 161.69324, 215.64265, 17.115429, 18.808159, 11.605783, 1.464602, 23.765022, 27.333698, 5.9699073, 0.38317743, 0.35822636, 7.4555554}
FF =
  {500.0, 200.0, 100.0, 1200.0, 100.0, 100.0, 100.0, 100.0, 2400.0, 200.0, 1800.0, 200.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 400.0, 200.0, 100.0, 100.0, 200.0, 300.0, 100.0, 100.0, 100.0, 200.0, 100.0, 100.0, 200.0, 700.0, 200.0, 600.0, 100.0, 100.0, 100.0, 2800.0, 100.0, 100.0, 100.0, 1000.0, 600.0, 100.0, 100.0, 600.0, 1000.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 100.0, 1400.0, 200.0, 100.0, 7300.0, 500.0, 100.0, 100.0, 100.0, 100.0, 100.0, 1700.0, 100.0, 200.0, 200.0, 100.0, 100.0, 100.0, 500.0, 100.0, 500.0, 2700.0, 200.0, 200.0, 200.0, 1200.0, 100.0, 2400.0, 100.0, 200.0, 100.0, 300.0, 100.0, 100.0, 100.0, 3300.0, 4600.0, 200.0, 400.0, 200.0, 400.0, 3800.0, 500.0, 1100.0, 100.0, 200.0, 1000.0, 600.0, 200.0, 100.0, 100.0, 100.0}
FA =
  {1.0, 2.0, 3.0, 4.0, 5.0, 6.0, 7.0, 8.0, 9.0, 10.0, 11.0, 12.0, 13.0, 14.0, 15.0, 16.0, 17.0, 18.0, 19.0, 20.0, 21.0, 22.0, 23.0, 24.0, 25.0, 26.0, 27.0, 28.0, 29.0, 30.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 39.0, 40.0, 41.0, 42.0, 43.0, 44.0, 45.0, 46.0, 47.0, 48.0, 49.0, 50.0, 51.0, 52.0, 53.0, 54.0, 55.0, 56.0, 57.0, 58.0, 59.0, 60.0, 61.0, 62.0, 63.0, 64.0, 65.0, 66.0, 67.0, 68.0, 69.0, 70.0, 71.0, 72.0, 73.0, 74.0, 75.0, 76.0, 77.0, 78.0, 79.0, 80.0, 81.0, 82.0, 83.0, 84.0, 85.0, 86.0, 87.0, 88.0, 89.0, 90.0, 91.0, 92.0, 93.0, 94.0, 95.0, 96.0, 97.0, 98.0, 99.0, 100.0, 101.0, 102.0, 103.0, 104.0, 105.0, 106.0, 107.0, 108.0, 109.0}
FGA =
  {0.0, 2.0, 4.0, 5.0, 8.0, 9.0, 10.0, 11.0, 12.0, 25.0, 27.0, 31.0, 32.0, 33.0, 34.0, 35.0, 36.0, 37.0, 38.0, 40.0, 41.0, 42.0, 43.0, 45.0, 47.0, 48.0, 49.0, 50.0, 51.0, 52.0, 53.0, 54.0, 59.0, 60.0, 61.0, 62.0, 63.0, 64.0, 72.0, 73.0, 74.0, 75.0, 78.0, 81.0, 82.0, 83.0, 87.0, 90.0, 91.0, 92.0, 93.0, 94.0, 95.0, 96.0, 97.0, 98.0, 99.0, 100.0, 101.0, 104.0, 105.0, 106.0, 118.0, 121.0, 122.0, 123.0, 124.0, 125.0, 126.0, 129.0, 130.0, 131.0, 132.0, 133.0, 134.0, 135.0, 137.0, 138.0, 141.0, 145.0, 147.0, 148.0, 150.0, 151.0, 152.0, 162.0, 163.0, 165.0, 166.0, 167.0, 168.0, 169.0, 170.0, 182.0, 193.0, 194.0, 196.0, 197.0, 198.0, 212.0, 215.0, 218.0, 219.0, 221.0, 225.0, 228.0, 230.0, 231.0, 232.0}
FGC =
  {2.0, 2.0, 1.0, 3.0, 1.0, 1.0, 1.0, 1.0, 13.0, 2.0, 4.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 2.0, 1.0, 1.0, 1.0, 2.0, 2.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 5.0, 1.0, 1.0, 1.0, 1.0, 1.0, 8.0, 1.0, 1.0, 1.0, 3.0, 3.0, 1.0, 1.0, 4.0, 3.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 3.0, 1.0, 1.0, 12.0, 3.0, 1.0, 1.0, 1.0, 1.0, 1.0, 3.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 2.0, 1.0, 3.0, 4.0, 2.0, 1.0, 2.0, 1.0, 1.0, 10.0, 1.0, 2.0, 1.0, 1.0, 1.0, 1.0, 1.0, 12.0, 11.0, 1.0, 2.0, 1.0, 1.0, 14.0, 3.0, 3.0, 1.0, 2.0, 4.0, 3.0, 2.0, 1.0, 1.0, 1.0}
FEA =
  {5.0, 2.0, 1.0, 12.0, 1.0, 1.0, 1.0, 1.0, 24.0, 2.0, 18.0, 2.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 4.0, 2.0, 1.0, 1.0, 2.0, 3.0, 1.0, 1.0, 1.0, 2.0, 1.0, 1.0, 2.0, 7.0, 2.0, 6.0, 1.0, 1.0, 1.0, 28.0, 1.0, 1.0, 1.0, 10.0, 6.0, 1.0, 1.0, 6.0, 10.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 1.0, 14.0, 2.0, 1.0, 73.0, 5.0, 1.0, 1.0, 1.0, 1.0, 1.0, 17.0, 1.0, 2.0, 2.0, 1.0, 1.0, 1.0, 5.0, 1.0, 5.0, 27.0, 2.0, 2.0, 2.0, 12.0, 1.0, 24.0, 1.0, 2.0, 1.0, 3.0, 1.0, 1.0, 1.0, 33.0, 46.0, 2.0, 4.0, 2.0, 4.0, 38.0, 5.0, 11.0, 1.0, 2.0, 10.0, 6.0, 2.0, 1.0, 1.0, 1.0}
DQF =
  {0, 0, 1, 0, 1, 1, 1, 1, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 0, 1, 1, 1, 0, 0, 1, 1, 1, 1, 1, 1, 1, 0, 1, 1, 1, 1, 1, 0, 1, 1, 1, 0, 0, 1, 1, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 1, 1, 0, 0, 1, 1, 1, 1, 1, 0, 1, 1, 1, 1, 1, 1, 0, 1, 0, 0, 0, 1, 0, 1, 1, 0, 1, 0, 1, 1, 1, 1, 1, 0, 0, 1, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 1, 1, 1}
nominal_satellite_subpoint_lat =
  {0.0}
nominal_satellite_subpoint_lon =
  {0.0}
nominal_satellite_height =
  {0.0}
geospatial_lat_lon_extent =
  {0.0}
OBIType =
  {0}
processing_parm_version_container =
  {0}
algorithm_product_version_container =
  {0}
}
